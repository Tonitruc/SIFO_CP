// megafunction wizard: %LPM_MUX%VBB%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: lpm_mux 

// ============================================================
// File Name: lpm_mux12.v
// Megafunction Name(s):
// 			lpm_mux
//
// Simulation Library Files(s):
// 			lpm
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 9.1 Build 350 03/24/2010 SP 2 SJ Web Edition
// ************************************************************

//Copyright (C) 1991-2010 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.

module lpm_mux12 (
	data0x,
	data10x,
	data11x,
	data1x,
	data2x,
	data3x,
	data4x,
	data5x,
	data6x,
	data7x,
	data8x,
	data9x,
	sel,
	result);

	input	[14:0]  data0x;
	input	[14:0]  data10x;
	input	[14:0]  data11x;
	input	[14:0]  data1x;
	input	[14:0]  data2x;
	input	[14:0]  data3x;
	input	[14:0]  data4x;
	input	[14:0]  data5x;
	input	[14:0]  data6x;
	input	[14:0]  data7x;
	input	[14:0]  data8x;
	input	[14:0]  data9x;
	input	[3:0]  sel;
	output	[14:0]  result;

endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Stratix II"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: CONSTANT: LPM_SIZE NUMERIC "12"
// Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_MUX"
// Retrieval info: CONSTANT: LPM_WIDTH NUMERIC "15"
// Retrieval info: CONSTANT: LPM_WIDTHS NUMERIC "4"
// Retrieval info: USED_PORT: data0x 0 0 15 0 INPUT NODEFVAL data0x[14..0]
// Retrieval info: USED_PORT: data10x 0 0 15 0 INPUT NODEFVAL data10x[14..0]
// Retrieval info: USED_PORT: data11x 0 0 15 0 INPUT NODEFVAL data11x[14..0]
// Retrieval info: USED_PORT: data1x 0 0 15 0 INPUT NODEFVAL data1x[14..0]
// Retrieval info: USED_PORT: data2x 0 0 15 0 INPUT NODEFVAL data2x[14..0]
// Retrieval info: USED_PORT: data3x 0 0 15 0 INPUT NODEFVAL data3x[14..0]
// Retrieval info: USED_PORT: data4x 0 0 15 0 INPUT NODEFVAL data4x[14..0]
// Retrieval info: USED_PORT: data5x 0 0 15 0 INPUT NODEFVAL data5x[14..0]
// Retrieval info: USED_PORT: data6x 0 0 15 0 INPUT NODEFVAL data6x[14..0]
// Retrieval info: USED_PORT: data7x 0 0 15 0 INPUT NODEFVAL data7x[14..0]
// Retrieval info: USED_PORT: data8x 0 0 15 0 INPUT NODEFVAL data8x[14..0]
// Retrieval info: USED_PORT: data9x 0 0 15 0 INPUT NODEFVAL data9x[14..0]
// Retrieval info: USED_PORT: result 0 0 15 0 OUTPUT NODEFVAL result[14..0]
// Retrieval info: USED_PORT: sel 0 0 4 0 INPUT NODEFVAL sel[3..0]
// Retrieval info: CONNECT: result 0 0 15 0 @result 0 0 15 0
// Retrieval info: CONNECT: @data 0 0 15 165 data11x 0 0 15 0
// Retrieval info: CONNECT: @data 0 0 15 150 data10x 0 0 15 0
// Retrieval info: CONNECT: @data 0 0 15 135 data9x 0 0 15 0
// Retrieval info: CONNECT: @data 0 0 15 120 data8x 0 0 15 0
// Retrieval info: CONNECT: @data 0 0 15 105 data7x 0 0 15 0
// Retrieval info: CONNECT: @data 0 0 15 90 data6x 0 0 15 0
// Retrieval info: CONNECT: @data 0 0 15 75 data5x 0 0 15 0
// Retrieval info: CONNECT: @data 0 0 15 60 data4x 0 0 15 0
// Retrieval info: CONNECT: @data 0 0 15 45 data3x 0 0 15 0
// Retrieval info: CONNECT: @data 0 0 15 30 data2x 0 0 15 0
// Retrieval info: CONNECT: @data 0 0 15 15 data1x 0 0 15 0
// Retrieval info: CONNECT: @data 0 0 15 0 data0x 0 0 15 0
// Retrieval info: CONNECT: @sel 0 0 4 0 sel 0 0 4 0
// Retrieval info: LIBRARY: lpm lpm.lpm_components.all
// Retrieval info: GEN_FILE: TYPE_NORMAL lpm_mux12.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL lpm_mux12.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL lpm_mux12.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL lpm_mux12.bsf TRUE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL lpm_mux12_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL lpm_mux12_bb.v TRUE
// Retrieval info: LIB_FILE: lpm
